
// @file add4.v
// @breif 4ビット加算器
// @author Yusuke Matsunaga (松永 裕介)
//
// Copyright (C) 2019 Yusuke Matsunaga
// All rights reserved.
//
// [概要]
// キャリー入力，キャリー出力つき4ビット加算器
//
// [入出力]
// a, b:   4ビット入力
// cin:    キャリー入力
// s:      4ビット出力
// cout:   キャリー出力
module add4(input [3:0]  a, b,
	    input 	 cin,
	    output [3:0] s,
	    output 	 cout);

endmodule // add4
